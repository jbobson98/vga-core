module vga_sync_generator #(

    // Horizontal pixel parameters (pixels)
    parameter HORZ_PIXELS = 640,
    parameter HORZ_FRONT_PORCH = 16,
    parameter HORZ_BACK_PORCH = 48,
    parameter HORZ_SYNC = 96,

    // Vertical pixel parameters (lines, 1 line is 1 pixel tall)
    parameter VERT_PIXELS = 480,
    parameter VERT_FRONT_PORCH = 10,
    parameter VERT_BACK_PORCH = 33,
    parameter VERT_SYNC = 2,

    // Width and height calculations
    parameter TOTAL_WIDTH = HORZ_PIXELS + HORZ_FRONT_PORCH + HORZ_BACK_PORCH + HORZ_SYNC,
    parameter WIDTH_BITS = $clog2(TOTAL_WIDTH + 1),
    parameter TOTAL_HEIGHT = VERT_PIXELS + VERT_FRONT_PORCH + VERT_BACK_PORCH + VERT_SYNC,
    parameter HEIGHT_BITS = $clog2(TOTAL_HEIGHT + 1)
    
)(
    input wire clk,
    input wire rst,
    output reg hsync,  // marks the beginning of a new line (generated by counting pixel clocks)
    output reg vsync,  // marks the beginning of a new data frame (generated by counting hsync transistions)
    output reg video_active,
    output wire [WIDTH_BITS-1 : 0] x_loc, // x coordinate of current pixel
    output wire [HEIGHT_BITS-1 : 0] y_loc  // y coordinate of current pixel
);


// Sync pulse reference points
localparam integer HORZ_SYNC_START = HORZ_PIXELS + HORZ_BACK_PORCH - 1;
localparam integer HORZ_SYNC_END = HORZ_PIXELS + HORZ_BACK_PORCH + HORZ_SYNC - 1;
localparam integer VERT_SYNC_START = VERT_PIXELS + VERT_FRONT_PORCH - 1;
localparam integer VERT_SYNC_END = VERT_PIXELS + VERT_FRONT_PORCH + VERT_SYNC - 1;

// Counters for tracking current pixel coordinate
wire x_loc_max;
flex_counter #(.MAX_COUNT(TOTAL_WIDTH-1), .WIDTH(WIDTH_BITS)) horizontal_counter 
    (.clk(clk), .rst(rst), .cen(1'b1), .maxcnt(x_loc_max), .count(x_loc));

wire y_loc_max;
flex_counter #(.MAX_COUNT(TOTAL_HEIGHT-1), .WIDTH(HEIGHT_BITS)) vertical_counter 
    (.clk(x_loc_max), .rst(rst), .cen(1'b1), .maxcnt(y_loc_max), .count(y_loc));

// Lines of each frame transmitted in order from top to bottom
// Pixels in each line are transmitted from left to right

// Line:  [ Active_Video  Front_Porch  H_Sync_Pulse  Back_Porch ]
// Frame: [ Active_Video(lines) Front_Porch V_Sync_Pulse Back_Porch ]
// HSYNC and VSYNC active low

// (i.e. the values lead genoration of syncpulse by 1 clock cycle)
// when horz_cnt = 655, hsync <= 1'b0; (HORZ_SYNC_START)
// when horz_cnt = 751, hsycn <= 1'b1;
// same for vsync at 489 and 491

always @(posedge clk or posedge rst) begin
    if(rst) begin
        hsync <= 1'b1;
        vsync <= 1'b1;
        video_active <= 1'b0;
    end else begin

        // Set video_active high only when we are in the active display region
        if((x_loc >= 0) && (x_loc < HORZ_PIXELS) && (y_loc >= 0) && (y_loc < VERT_PIXELS)) begin
            video_active <= 1'b1;
        end else begin
            video_active <= 1'b0;
        end

        // Set hsync pulse
        if((x_loc >= HORZ_SYNC_START) && (x_loc <= HORZ_SYNC_END)) begin
            hsync <= 1'b0;
        end else begin
            hsync <= 1'b1;
        end

        // Set vsync pulse
        if((y_loc >= VERT_SYNC_START) && (y_loc <= VERT_SYNC_END)) begin
            vsync <= 1'b0;
        end else begin
            vsync <= 1'b1;
        end

    end
end

endmodule