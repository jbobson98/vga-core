// Top level module for VGA experimentation on the Digilent BASYS 3 development board

module vga_core (
    input wire clk,
    input wire rst,
    output wire hsync,
    output wire vsync,
    output wire [3:0] red,
    output wire [3:0] green,
    output wire [3:0] blue
);

// Instantiate 25MGHZ clock


// Debounce reset


// instantiate vga_sync_gen



endmodule