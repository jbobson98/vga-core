module resolution_selector (
    // clk input, rst, mux select
    // ooutput regs
    intput wire clk,
    input wire rst,
    input wire [3:0] sel,


);









    // HORZ_PIXELS = 11bits
    // VERT_PIXELS = 11bits
    // 2^9 for each porch and pulse





    // all at 60hz
    // 640x480 #
    // 800x600 #
    // 1024x768 #
    // 1280x720 #
    // 1280x1024 #
    // 1600x1200 #
    // 1920x1080 #




endmodule